module shift_ram 
  (
   clk,
   ce,
   d,
   q
   );

   input          clk;
   input 		  ce;
   input [7 : 0]  d;
   output [7 : 0] q;
   
endmodule
