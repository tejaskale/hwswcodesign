library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-------------------------------------------------------------------------------

entity pipe_control_logic is
  port (i_empty : in  std_logic;
        o_full  : in  std_logic;
        enable  : out std_logic);
end pipe_control_logic;

-------------------------------------------------------------------------------

architecture behavioral of pipe_control_logic is

begin

-- 
-- WRITE YOUR CODE HERE
--

end behavioral;

